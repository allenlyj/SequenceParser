`timescale 1ns/1ps
`include "parser.sv"
module tb_parser;

    //Input signals
    reg clk = 0, reset = 1'b1, dataInVal = 0, dataOutReady = 0, dataInLast = 0;
    reg [31:0] dataIn = 0;
    //Output signals
    wire dataInReady, dataOutVal, packetLost;
    wire [0:295] dataOut;
    parser yaojie(.clk(clk), .reset_b(reset), 
                   .dataIn(dataIn), .dataIn_val(dataInVal), 
                   .dataIn_ready(dataInReady), .dataIN_last(dataInLast),
                   .dataOut(dataOut), .dataOut_val(dataOutVal),
                   .dataOut_ready(dataOutReady), .packetLost(packetLost));
    

    always begin
        clk = 1'b0;
        #5;
        clk = 1'b1;
        #5;
    end

    task sendPacket(input int stream, input int seq, input int length) begin
        reg[15:0] streamLE = {stream[7:0], stream[15:8]};
        reg[31:0] seqLE = {seq[7:0], seq[15:8], seq[23:16], seq[31:24]};
        reg[15:0] lengthLE = {length[7:0], length[15:8]};
        int cycles = length/4;
        int i = 0;
        dataInVal = 1'b1;
        while (i < cycles) begin
            @ (posedge clk) begin
                if (i == 0)
                    dataIn = {lengthLE, streamLE};
                else if (i == 1)
                    dataIn = seqLE;
                else
                    dataIn = 32'h01234560 + i;
                if (dataInReady)
                    i = i + 1;
            end
        dataInVal = 1'b0;
    end

    initial begin
        $monitor("valid=%d last=%d data=%8x ready=%d", dataInVal, dataInLast, dataIn, dataInReady);
        reset = 1'b0;
        #50ns reset = 1'b1;
        sendPacket(12, 1, 20);
        sendPacket(13, 1, 25);
        sendPacket(12, 3, 39);
        #200 $finish;
    end
    always @ (posedge clk)
        $display ("T=%0t dataOut=0x%0h %x", $time, dataOut, yaojie.seqs[5]);
    always @ (negedge clk)
        $display ("T=%0t dataOut=0x%0h", $time, dataOut);
endmodule