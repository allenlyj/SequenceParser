module parser(clk, reset_b, dataIn, dataIn_val, dataIn_ready, dataIn_last, //receive interface
               dataOut, dataOut_val, dataOut_ready, packetLost); //send interface
    
    input clk, reset_b, dataIn_val, dataIN_last, dataOut_ready;
    input [31:0] dataIn;
    output dataIn_ready, dataOut_val;
    output reg packetLost = 0;
    output [0:295] dataOut;

    reg [0:295] outputPrepare = 0;
    reg [0:295] outputFinal = 0;
    reg [31:0] seqs [0:31];
    reg outputPending = 0;
    localparam [1:0] IDLE = 0;
    localparam [1:0] GET_2ND_WORD = 1;
    localparam [1:0] GET_DATA = 2;
    localparam [1:0] COMMIT_OUTPUT = 3;
    reg [1:0] receiverState = IDLE;
    reg [15:0] bytesLeft = 0;
    reg [15:0] currentStream = 0;
    reg [31:0] currentSeq = 0;
    reg [3:0] currentOutputIndex = 0;
    wire canMoveForward;
    wire [31:0] maskedInput;
    wire sequenceValid;
    wire [4:0] currentStream;

    integer i;

    assign dataIn_ready = !(outputPending or receiverState == COMMIT_OUTPUT);
    assign dataOut_val = outputPending;
    assign canMoveForward = !outputPending & dataIn_val;
    assign currentSeqTrimmed = currentSeq[4:0];
    assign sequenceValid = (currentSeq == seqs[currentSeqTrimmed] + 1);

    always @ (*) begin
        if (!dataIn_last) 
            maskedInput = dataIn;
        else begin
            case (bytesLeft)
                1 : maskedInput = {dataIn[31:24], 24'd0};
                2 : maskedInput = {dataIn[31:16], 16'd0};
                3 : maskedInput = {dataIn[31:8], 8'd'0};
                4 : maskedInput = 
                default : maskedInput = 0; //Bad format, should not happen or should trigger error flag

            endcase
        end
    end

    always @ (posedge clk)
        if (!reset_b) begin
            outputPending <= 0;
            for (i = 0; i <= 31; i = i+1) begin
                seqs[i] <= 0;
            end
            receiverState <= IDLE;
            outputPrepare <= 0;
        end else begin
            // Only move forward if there is incoming data and no pending transaction
            case(receiverState)
            IDLE:
                if (canMoveForward) begin
                    bytesLeft <= dataIn[31:16]-4;
                    currentStream <= dataIn[15:0];
                    receiverState <= GET_2ND_WORD;
                end
            GET_2ND_WORD:
                if (canMoveFoward) begin
                    bytesLeft <= bytesLeft - 4;
                    currentSeq <= dataIn;
                    receiverState <= GET_DATA;
                    currentOutputIndex <= 0;
                end
            GET_DATA:
                if (canMoveFoward) begin
                    outputPrepare[currentOutputIndex*32 : currentOutputIndex:32+31] <= maskedInput;
                    currentOutputIndex <= currentOutputIndex + 1;
                    bytesLeft <= bytesLeft - 4;
                    if (dataIn_last) begin
                        receiverState <= COMMIT_OUTPUT;
                        packetLost <= !sequenceValid
                        seqs[currentSeqTrimmed]
                    end

                end
            endcase
        end



        
endmodule